CMOS Buffer
vdd 4 0 dc 5v
vina 2 0 pulse(0v 5v 0 1ns 1ns 10ns 20ns)

m1 2 1 4 4 pmod l=1u w=100u
m2 2 1 0 0 nmod l=1u w=40u
m3 3 2 4 4 pmod l=1u w=100u
m4 3 2 0 0 nmod l=1u w=40u

.model nmod nmos vto=1v kp=200u
.model pmod pmos vto=-v kp=80u

.tran 0.1ns 120ns
.control
run
plot v(5) v(2) v(1)
.endc
.end
