a simple circuit with 3 resistors in parallel
v1 1 0 dc 9v
r1 2 0 5k
r2 3 0 10k
r3 4 0 15k

vr1 1 2 dc 0
vr2 1 3 dc 0
vr3 1 4 dc 0

.dc v1 9 9 1
.print dc v(2,0) v(3,0) v(4,0)
.print dc i(vr1) i(vr2) i(vr3)
.plot 
.end
