a'b'+c'
vdd 7 0 dc 5v
vina 1 0 pulse(0V 5V 0 1ns 1ns 10ns 20ns)
vinb 2 0 pulse(0V 5V 0 1ns 1ns 15ns 20ns)
vinc 3 0 pulse(0V 5V 0 1ns 1ns 5ns 20ns)

*upper half
m1 6 1 7 7 mos1 l=1u w=100u
m2 5 2 6 6 mos1 l=1u w=100u
m3 5 3 7 7 mos1 l=1u w=100u

*lower half
m4 5 1 4 4 mos2 l=1u w=40u
m5 5 2 4 4 mos2 l=1u w=40u
m6 4 3 0 0 mos2 l=1u w=40u

.model mos2 nmos vto=1v kp=200u
.model mos1 pmos vto=-1v kp=80u

.tran 0.1ns 120ns
.control
run
plot v(5) v(1) v(2) v(3)
.endc
.end
