Logic Function ((a'+b')c') using CMOS logic
* ((a'+b')c') = a'c'+b'c'
vdd 7 0 dc 5v
*input voltage
vin1 1 0 pulse(0V 5V 0 1ns 1ns 10ns 20ns)
vin2 2 0 pulse(0V 5V 0 1ns 1ns 15ns 20ns)
vin3 3 0 pulse(0V 5V 0 1ns 1ns 5ns 20ns)

* upper half pmos
m1 6 1 7 7 mos1 l=1u w=100u
m2 6 2 7 7 mos1 l=1u w=100u
m3 5 3 6 6 mos1 l=1u w=100u

* lower half nmos
m4 5 2 4 4 mos2 l=1u w=40u
m5 4 1 0 0 mos2 l=1u w=40u
m6 5 3 0 0 mos2 l=1u w=40u

.model mos2 nmos vto=1v kp=200u
.model mos1 pmos vto=-1v kp=80u

.tran 0.1ns 120ns
.control
run
plot v(5) v(1) v(2) v(3)
.endc
.end
