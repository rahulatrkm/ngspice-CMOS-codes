CMOS transmission gate
vdd 4 0 dc 5v
vina 2 0 pulse(0v 5v 0 1ns 1ns 10ns 20ns)
vinb 1 0 pulse(0v 5v 0 1ns 1ns 5ns 20ns)
vinbbar 3 0 pulse(5v 0v 0 1ns 1ns 10ns 20ns)
m1 5 1 2 0 mos1 w=40u l=1u
m2 2 3 5 4 mos2 w=100u l=1u

.model mos1 nmos vto=1v kp=200u
.model mos2 pmos vto=-1v kp=80u

.tran 0.1ns 120ns
.control
run
plot v(5) v(2) v(1)
.endc
.end
