Tristate Inverter
vdd 7 0 dc 5v

*input voltages
vin1 1 0 pulse(0V 5V 0 1ns 1ns 10ns 20ns)
vin2 2 0 pulse(0V 5V 0 1ns 1ns 10ns 20ns)
vin2bar 3 0 pulse(5V 0V 0 1ns 1ns 10ns 20ns)

*upper half
m1 6 1 7 7 mos1 l=1u w=100u
m2 5 3 6 6 mos1 i=1u w=100u

*lower half
m3 5 2 4 4 mos2 l=1u w=40u
m4 4 1 0 0 mos2 l=1u w=40u

.model mos1 pmos vto=-1v kp=80u
.model mos2 nmos vto=1v kp=200u

.tran 0.1ns 120ns
.control
run
plot v(5) v(2)
