CMOS Buffer
vdd 4 0 dc 5v
vin1 1 0 pulse(0v 5v 0 1ns 1ns 10ns 20ns)

m1 2 1 4 4 mos2 l=1u w=100u
m2 2 1 0 0 mos1 l=1u w=40u
m3 3 2 4 4 mos2 l=1u w=100u
m4 3 2 0 0 mos1 l=1u w=40u

.model mos1 nmos vto=1v kp=200u
.model mos2 pmos vto=-1v kp=80u

.tran 0.1ns 120ns
.control
run
plot v(5) v(2) v(1)
.endc
.end
