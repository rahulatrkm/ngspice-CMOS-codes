.model MOSN NMOS
.model MOSP PMOS

