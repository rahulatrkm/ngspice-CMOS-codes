Logic Function ((a'+b')c') using CMOS logic
* ((a'+b')c') = a'c'+b'c'
vdd 8 0 dc 5v
* upper half pmos
m1 8 1 7 8 mos1 l=10u w=100u
.model mos1 pmos vto=1.5v kp=200u
m2 8 3 6 8 mos2 l=10u w=100u
.model mos2 pmos vto=1.5v kp=200u
m3 7 2 5 7 mos3 l=10u w=100u
.model mos3 pmos vto=1.5v kp=200u
m4 6 2 5 6 mos4 l=10u w=100u
.model mos4 pmos vto=1.5v kp=200u
* lower half nmos
m5 5 1 6 6 mos5 l=10u w=100u
.model mos5 nmos vto=1.5v kp=200u
m6 5 2 6 6 mos6 l=10u w=100u
.model mos6 nmos vto=1.5v kp=200u
m7 4 2 7 7 mos7 l=10u w=100u
.model mos7 nmos vto=1.5v kp=200u
m8 4 3 7 7 mos8 l=10u w=100u
.model mos8 nmos vto=1.5v kp=200u
vin1 1 0 pulse(2 5 0 0 0 100ns 800ns)
vin2 2 0 pulse(2 5 0 0 0 100ns 800ns)
vin3 3 0 pulse(2 5 0 0 0 100ns 800ns)
.tran 10ns 1200ns
.control
run
plot v(5) v(1) v(2) v(3)
.endc
.end
